// Simplest possible Verilog program to verify environment.
module main;
  initial 
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule